                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                                S02B0000433A5C55736572735C44616E5C417070446174615C4C6F63616C5C54656D705C61726475696E6F5F9D
S113040097410000938181E097440000938404ABFA
S113041017340000130484696F00C0002300040033
S113042013041400E31C94FE173400001304845CCA
S1130430973400009384445C138900006F0000012A
S11304400325040013044400E7000500E31A94FEA6
S10B0450930009006F00C000D5
S11304581385018A6F00903C130101FF2324810056
S1130468370400002326110013040400EF108073DE
S1130478EF008001EF004004E30E04FE9700000043
S1130488E780C0B76FF01FFF130101FF2324810029
S11304981385018A23261100EF10C04C1385018AA5
S11304A8EF1000281385018A032481008320C100EA
S11304B8130101016F100042130101FA232C810476
S11304C8232A91049384818A03A50400232E11040A
S11304D823282105232631052324410523225105F8
S11304E8232C8103232A910323206105232E7103DE
S11304F82328A1032326B103EF10406C93050500BC
S1130508EF10D07F930A050003A50400B707008005
S11305183345F500EF10806A93050500EF10107E4F
S11305282324A1001385018AEF10801F930C200057
S11305381384818A374A0000374C00003749000089
S1130548B749000013850C00EF20100AB7470000D4
S113055803A6078483A64784EF20102A130B0500FB
S113056803250400938B0500EF20406E13060B004F
S113057893860B00EF101032EF304011EF10006437
S1130588B747000083A507812320A10003250400A1
S1130598EF10D076EF20806B13060B0093860B00C8
S11305A8EF10502FEF30800EEF104061930B0500D1
S11305B813953C00EF20900C93850A00130D050059
S11305C8EF10D073232EA100EF204076B747000028
S11305D883A5478183270100931D050193DD0D4100
S11305E813850700EF209061B747000083A5878132
S11305F8130B0500938C1C00EF105070EF20007350
S1130608131E0501135E0E4113060E001307100096
S11306189306200093850D001385018A232CC101BC
S1130628EF00106C8325810013050D00EF10106D89
S1130638232AA100EF20806F83254981131D05011A
S113064813850B00EF20905B83A58981930B05002C
S1130658135D0D41EF10906AEF20406D13130501EF
S113066813530341130603009306200013071000D5
S113067893050D001385018A23286100EF00506655
S11306888325498113850B00EF105067EF20006A1A
S113069883254981131705011357074113050B00D7
S11306A82320E100EF109065EF2040680327010044
S11306B8131605019307100093060D0013560641FF
S11306C893850D001385018AEF00902013850C0093
S11306D8EF20807103260A8483264A84374B00005E
S11306E8EF2090112320A100032504002322B10048
S11306F8EF20C0550326010083264100EF1090190E
S1130708EF20D078EF10804B83254981EF20104FDC
S113071883A58981EF10905EEF204061032FC1010A
S11307288325CB81131705011357074113050F00C0
S11307382326E100EF10905CEF20405F032E810137
S11307480327C1009316050113060E009307100032
S113075893D6064193850D001385018AEF0050173F
S113076883250C8103250400EF105059EF20004E17
S11307780326010083264100EF10D011EF201071E9
S1130788EF10C04383254981EF20504783A5898111
S1130798EF10D056EF208059832E41018325CB8159
S11307A8131705011357074113850E002320E10091
S11307B8EF10D054EF2080570323010103270100D1
S11307C8931605019307100093D6064113060300F8
S11307D893050D001385018AEF00900F9307F0002D
S11307E8E392FCD603250400938B0189EF2000468D
S11307F81306000093060000EF10D009EF201069DB
S1130808B7490000839C0B00EF10403B83A5098285
S113081837490000930D2000EF20503E9305050052
S113082803254982EF209065EF2040509315050178
S1130838930710001307800093068000138601862F
S113084813850C0093D50541EF00106E03250400B1
S113085883AC0B00EF20803F03260A8483264A8456
S1130868938CAC00939C0C01EF10D002EF20106223
S1130878EF10C03483A5098293DC0C41EF201038B3
S11308889305050003254982EF20505FEF20004AB5
S11308989315050113078000930710009306800041
S11308A81386818513850C0093D50541EF00D06725
S11308B80325040003AA0B00EF204039B7470000C2
S11308C803A6878483A6C784130A4A01131A0A0154
S11308D8EF10407CEF20905BEF10402E83A5098237
S11308E8135A0A41EF2090319305050003254982E4
S11308F8EF20D058EF20804393150501130780009B
S113090813868186930710009306800013050A0056
S113091893D50541EF0050610325040003AA0B0099
S1130928EF20C032B747000003A6078583A6478592
S1130938130AEA01131A0A01EF10C075EF201055C3
S1130948EF10C02783A50982135A0A41EF20102B00
S11309589305050003254982EF205052EF20003DFE
S113096893150501130780001386818693071000E9
S11309789306800013050A0093D50541EF00D05A69
S11309880325040003AA0B00EF20402CB7470000FE
S113099803A6878583A6C785130A8A02131A0A0140
S11309A8EF10406FEF20904EEF10402183A509828D
S11309B8135A0A41EF209024930505000325498220
S11309C8EF20D04BEF2080369315050113078000E4
S11309D893071000930680001386018713050A0005
S11309E893D50541EF0050540325040003AA0B00D6
S11309F8EF20C025B747000003A6078683A64786CD
S1130A08130A2A03131A0A01EF10C068EF201048CA
S1130A18EF10C01A83A50982135A0A41EF20101E49
S1130A289305050003254982EF205045EF20003047
S1130A38931505011307800093071000930680009F
S1130A481386818313050A0093D50541EF00D04D21
S1130A580325040003AA0B00EF20401FB74700003A
S1130A6803A6878683A6C786130ACA03131A0A012C
S1130A78EF104062EF209041EF10401483A50982E3
S1130A88135A0A41EF20901793050500032549825C
S1130A98EF20D03EEF20802993150501130780002D
S1130AA893071000930680001386018413050A0037
S1130AB893D50541EF0050470325040003AA0B0012
S1130AC8EF20C018B747000003A6078783A6478707
S1130AD8130A6A04131A0A01EF10C05BEF20103BD3
S1130AE8EF10C00D83A50982135A0A41EF20101193
S1130AF89305050003254982EF205038EF20002391
S1130B0893150501130780009307100093068000CE
S1130B181386818713050A0093D50541EF00D04059
S1130B280325040003AA0B00EF204012B747000076
S1130B3803A6878783A6C787130A0A05131A0A0117
S1130B48EF104055EF209034EF10400783A5098239
S1130B58135A0A41EF20900A930505000325498298
S1130B68EF20D031EF20801C931505011307800076
S1130B7893071000930680001386018513050A0065
S1130B8893D50541EF00503A0325040003AA0B004E
S1130B98EF20C00BB747000003A6078883A6478841
S1130BA8130AAA05131A0A01EF10C04EEF20102EDB
S1130BB8EF10C00083A50982135A0A41EF201004DC
S1130BC89305050003254982EF20502BEF200016DA
S1130BD893150501130780009307100093068000FE
S1130BE81386018813050A0093D50541EF00D03315
S1130BF80325040003AA0B00EF204005B7470000B3
S1130C0803A6878883A6C788130A4A06131A0A0103
S1130C18EF104048EF209027EF00507A83A509820F
S1130C28135A0A41EF20807D930505000325498264
S1130C38EF20D024EF20800F9315050113078000BF
S1130C4893071000930680001386818413050A0015
S1130C5893D50541EF00502D0325040003AA0B008A
S1130C68EF10D07EB747000003A6078983A64789FB
S1130C78130AEA06131A0A01EF10C041EF201021E3
S1130C88EF00D07383A50982135A0A41EF20007735
S1130C989305050003254982EF20501EEF20000923
S1130CA8931505011307800093071000930680002D
S1130CB81386018713050A0093D50541EF00D02652
S1130CC80325040003AA0B00B74B0000EF101078AB
S1130CD8B747000003A6878983A6C789130A8A072A
S1130CE8131A0A01EF10003BEF20501AEF00106DA1
S1130CF883A50982135A0A41B7490000EF200070FE
S1130D089305050003254982EF205017EF200002C0
S1130D1893150501930710001307800093068000BC
S1130D281386818893D5054113050A00EF00D01F67
S1130D38B747000083A5878213850A00EF20006C5B
S1130D4893880189130D0500374C00009305600052
S1130D5813850D0023281101EF10C022EF20001283
S1130D681309050013850D00EF200008B74700009C
S1130D7803A6078A83A6478A938D1D00EF20C02700
S1130D88130A050003250400938A0500EF10106C6C
S1130D9893860A0013060A00EF10C02FEF20100FE5
S1130DA8EF00D061B747000083A5C782930C050004
S1130DB813050D00EF108074EF10507E8325CB814E
S1130DC81377F50F13850C002324E100EF2000634B
S1130DD8B747000083A50783EF104072EF10107522
S1130DE8131605011356064193050D001305090052
S1130DF82320C100EF108070EF1050730327810087
S1130E08032601009315050193064000930710007B
S1130E1893D505411385018AEF00D001B747000037
S1130E2883A5478303250400EF10406DEF00105994
S1130E38930C050083254C8303250400EF10006CF4
S1130E48EF10D06013060A0093860A00EF1080247E
S1130E58EF20D003EF00905683254C832320A10074
S1130E6803250400EF108069EF00505583A5CB8259
S1130E78EF10C068EF109072832601008325CB81A0
S1130E881377F50F138506002324E100EF2000579C
S1130E9883A50983EF108066EF10506913160501C6
S1130EA81356064193850C00130509002320C1003D
S1130EB8EF10C064EF109067032781000326010038
S1130EC893150501930710009306400093D5054137
S1130ED81385018AEF000076B74C000083A58C8344
S1130EE803250400EF108061EF00504D83A58C8327
S1130EF82326A10003250400EF104060EF101055CD
S1130F0893860A0013060A00EF10C018EF20007831
S1130F18EF00D04A83A58C83130A05000325040037
S1130F28EF10C05DEF00904983A5CB82EF10005D00
S1130F38EF10D0668325CB811377F50F13050A00CC
S1130F482324E100EF20804B83A50983EF10005B85
S1130F58EF10D05D0323C100131605011356064193
S1130F6893050300130509002320C100EF1000595D
S1130F78EF10D05B032781000326010093150501B8
S1130F88930710009306400093D505411385018A01
S1130F98EF00406A9307400183280101E398FDDAD2
S1130FA883A708001307E0F79387F7FF6384E7062E
S1130FB80325040023A0F800EF105049B7470000A8
S1130FC803A6078A83A6478AEF10C00CEF20006C9B
S1130FD82320A400032481058320C10503290105D6
S1130FE88329C104032A8104832A4104032B0104AD
S1130FF8832BC103032C8103832C4103032D010399
S1131008832DC1021385018A832441051301010636
S11310186F00500C930710086FF09FF9130101FF3C
S1131028232611002324810013040500EF009016E1
S1131038930700012311F40023020400130500019F
S1131048EF0090158320C10023100400230304003B
S113105803248100130101016780000013150501B1
S1131068135505019307F00763ECA704939505014D
S113107893D505019307F00363E4B70413F77500E8
S113108893F5850F9395450093071000B305B500B4
S1131098B397E700939505019386018B93D50501D2
S11310A8B386B60093F7F70F83C606001387018B40
S11310B8630A0600B3E7F600B305B7002380F5001A
S11310C86780000093C7F7FFB3F7F6006FF0DFFE01
S11310D8130101FD232C4101330AC7402324810154
S11310E8138C07009357FA4133CA4701232A510145
S11310F8B38AB640330AFA4093D7FA41B3CA5701C0
S11311082324810223229102232E31012326110252
S1131118232021032328610123267101232291011D
S1131128B38AFA40138405009304060093890600E1
S113113863DA4A01930907001304060013870600BB
S11311489384050063DE89009387040093040700F1
S11311581387070093070400138409009389070081
S1131168330B9740B38B89409357FB41939B0B01F7
S113117833CB670193DB0B01330BFB4093970B01D4
S113118893D7074113D9F7013309F90013591940C3
S1131198930C100063C4E400930CF0FF63C2890647
S11311A813060C0063D84A0593050400138504004C
S11311B833096941EFF09FEA9317090193D70701AF
S11311C81399070113590941635E0900B3849C000C
S11311D83389FB00939404011319090193D404413E
S11311E8135909411304140013140401135404413A
S11311F86FF0DFFA93850400130504006FF05FFBBA
S11312088320C102032481028324410203290102A9
S11312188329C101032A8101832A4101032B010186
S1131228832BC100032C8100832C4100130101038B
S113123867800000130101FD232481022322910207
S11312482320210323261102232E310113890500AB
S1131258B304D60013040000634406001304060014
S113126813140401135404419309000493870400DC
S113127863D49900930700046354F402931504019A
S11312881306070093D50541130509002326E10039
S1131298EFF0DFDC130414000327C1006FF01FFD17
S11312A88320C10203248102832441020329010209
S11312B88329C1011301010367800000130101FBA5
S11312C823286103130B050013950601232E31030C
S11312D8232C410313550501138A050093091000B3
S11312E89305E0FF2324810423202105232A5103A5
S11312F813890700232671032324810323229103DE
S1131308130C07002320A103930A06001384060084
S11313182326110423229104232EB101930B0800E0
S1131328B389A940EF00104693771C00931C05016C
S113133813140401131A0A01939A0A0113091900D0
S113134893DC0C4113540441130D00002324F100D1
S1131358135A0A0193DA0A011379F90F137C2C0042
S113136863528D1463C80902938C2C0093970C0163
S113137893D707011304F4FFB38937011314040145
S1131388939C0701939909011354044193DC0C417C
S113139893D9094193041D009394040193D404013F
S11313A8939D140093871D00B38937018327810017
S11313B8139D040193990901135D0D4193D90941C2
S11313C8638807069317040193D707013386FA4005
S11313D893161400B3059A00B306D9001316060130
S11313E89395050113870B0093F6F60F13560641E0
S11313F893D5054113050B002326F100EFF09FE375
S11314088327C10033869A40B306B901B305FA00AD
S1131418131606019395050113870B0093F6F60F2F
S11314281356064193D5054113050B00EFF09FE0D1
S1131438E3080CF29317040193D707013386FA40A3
S113144893161400B3059A40B306D900131606017F
S11314589395050113870B0013050B0093F6F60FFC
S11314681356064193D505412326F100EFF09FDC7E
S11314788327C10033869A40B306B901B305FA40FD
S1131488131606019395050113870B0093F6F60FBF
S11314981356064193D5054113050B00EFF09FD968
S11314A86FF01FEC8320C1040324810483244104C6
S11314B8032901048329C103032A8103832A4103DD
S11314C8032B0103832BC102032C8102832C4102C9
S11314D8032D0102832DC10113010105678000005A
S11314E8130101FD2324810213840600232291029F
S11314F893961600930406003306864093861600D6
S11315081316060193F6F60F1356064123202103FA
S1131518232E31012326110213090500938905009E
S11315282326E100EFF01FD193060400032481026F
S11315380328C1008320C10213860400938509008F
S1131548832441028329C1011305090003290102E7
S11315589307000013073000130101036FF01FD62F
S113156813150601135505019307F00363E2A70C4D
S1131578B386B6001398060113580841635A000B42
S11315889307F00763C6B70A9387050063D4050079
S113159893070000939507019307000893D5054125
S11315A89306080063D407019306000813563640CF
S11315B8931776003386B7009387018BB386B640BA
S11315C8B387C70093051000137675003396C500DA
S11315D893F6F60F1376F60F63060702631AB70439
S11315E89305F00F9386F6FF93F6F60F6382B6041D
S11315F803C70700938717003367E600A38FE7FE46
S11316086FF05FFE1346F6FF1376F60F9305F00F9F
S11316189386F6FF93F6F60F638CB60003C70700AC
S1131628938717003377E600A38FE7FE6FF05FFE1A
S113163867800000130101FE23244101130A0700F7
S113164813870700232E1100232C8100232A9100DD
S113165823282101232631012322510193840700E1
S11316689309060013090500938A050013840600EC
S1131678EFF01FEF1306FAFF3306360113160601BF
S1131688138704009306040093850A0013050900D0
S113169813560641EFF0DFEC1387040093060A00A3
S11316A81386090093850A0013050900EFF09FB813
S11316B89305F4FF03248101B38555018320C101F7
S11316C8832A41001387040093060A0083244101F6
S11316D8032A810013860900130509008329C10020
S11316E8032901019395050193D5054113010102CD
S11316F86FF05FB4B335B000B305B04093F5F50FA0
S1131708930700001387018B930600403306F70004
S11317182300B60093871700E39AD7FE678000007A
S1131728930500006FF01FFD3308D50063420818C5
S11317381308F007634EA8163308B700634A08165F
S11317481308F0036346B81613D8F541B348B80034
S1131758130101FFB3880841137878003308B800EF
S113176823268100232491002322210123203101EF
S113177893F878001358384063D80500930580001F
S11317881308F8FFB3881541935E37001377770081
S113179863040700938E1E0013137800B305A30097
S11317A81383018B130F8000130708003303B3005E
S11317B8B38E0E01930FF0FF1304F007B3041F4117
S11317C893021000130970006388EE0C6306E70D9A
S11317D86348F70B130E0000930303086352DE0AF1
S11317E8B305AE00634EB40863C005066302F70B85
S11317F83308C60103480800B309C30183850900F7
S11318083318180113188801135888416392570430
S1131818B3E505012380B90063880802630627033A
S11318283308C60103480800B389C3018385090046
S113183833589840131888011358884163965702FF
S1131848B3E505012380B900130E1E006FF01FF9DC
S1131858639807001348F8FFB3F505016FF09FFB81
S1131868B3C505016FF01FFB639807001348F8FF21
S1131878B3F505016FF01FFDB3C505016FF09FFCBB
S113188813071700130303083306D6006FF0DFF3BA
S1131898E39808F86FF05FFB0324C10083248100F8
S11318A80329410083290100130101016780000015
S11318B86780000037460000930505009307100071
S11318C813070001930680051306868A1305400151
S11318D86FF09FE5930500001385018B6F00C0131B
S11318E8130101FE232C8100232A910023282101BE
S11318F823263101232E1100930405009389050042
S1131908130400FF1309900113850400EFF05FE14D
S113191813050400E7800900138504001304140068
S1131928EFF05FFB131404011305F0001354044192
S1131938EF000018E31A24FD032481018320C10168
S113194883244101032901018329C10013050019D6
S1131958130101026F00C015B72500009385C58BDC
S11319686FF01FF8130101FF2326110023248100BF
S113197813040500EF00000A13050400EFF09FF5B7
S113198813050400032481008320C100130101010D
S11319986FF09FFC678000002386A18A678000009F
S11319A8130101FF23248100130400F18327040099
S11319B83717F040130707A023261100B3F7E700F1
S11319C82320F40083270400370710001307072097
S11319D8B3E7E7002320F400832704003707F0FF68
S11319E81307F7DFB3F7E7002320F400930510008B
S11319F81305D000EF00000F832704008320C100E3
S1131A0893E707402320F400032481001301010114
S1131A18678000006FF0DFF8832700F13707800044
S1131A283716F0FFB3E7E700B706C0FF2328F0F046
S1131A38930805401306F6FF9386F6FF370840001F
S1131A48032700F13377C7002328E0F08347050014
S1131A58638A0700032700F19397C700B3E7E700F9
S1131A682328F0F06384050023000500032700F110
S1131A78130515003377D7002328E0F0032700F176
S1131A88336707012328E0F0E31C15FB032700F163
S1131A98B70640FF9386F6FF3377D7002328E0F094
S1131AA8832700F1B3E707012328F0F067800000DB
S1131AB86F004000F32710C0378701001306F0FFBA
S1131AC81307076A1305F5FF6314C5006780000050
S1131AD8B387E700F32610C0B386D740E34CD0FEA3
S1131AE86FF05FFE83A74189637CF50AB74700005E
S1131AF893878795131515003305F500834705006B
S1131B08374700001307479F93F7770093972700F9
S1131B18B387E70003A70700930700806312F70859
S1131B28930710006382F506638C05029306200070
S1131B386398D5060346050083254080135636006E
S1131B48B397C70093C6F7FFB3F6B6002322D08035
S1131B5883260700B3E7D7002320F7006780000037
S1131B68034605008326408013563600B397C70002
S1131B7893C7F7FFB3F6F6002322D0808326070025
S1131B88B3F7D7006FF05FFD834705000327408054
S1131B9893D73700B395F500B3E5E5002322B08069
S1131BA86780000023260080232A00809307F0FF23
S1131BB82324F0802328F08067800000B7470000C2
S1131BC883A587A3130101FE232E1100232C810072
S1131BD8232A910023282101B7440000232441012A
S1131BE8232251012326310197020000E780822035
S1131BF81304050097120000E780820503A684A059
S1131C0883A6C4A0130A0500938A0500971200004E
S1131C18E78042CD1389040063460502B7400000FB
S1131C2803A600A183A640A113050A0093850A0010
S1131C3897220000E78002A397220000E78042A5CC
S1131C4813040500B74400001305040097120000AC
S1131C58E780020003A684A183A6C4A19309050012
S1131C68138A050097120000E78002D16356050223
S1131C78B742000003A602A183A642A11385090066
S1131C8893050A0097020000E780024197220000AA
S1131C98E78002A01304050013050400971200004E
S1131CA8E78002FB37430000032603A2832643A2EE
S1131CB893090500938A050097120000E78082C201
S1131CC863440502032589A08325C9A01386090056
S1131CD893860A0097220000E780C29897220000A2
S1131CE8E780029B13040500130504009712000003
S1131CF8E78002F6B743000003A683A283A6C3A223
S1131D0813090500138A050097120000E780C2C66C
S1131D186354050203A584A183A5C4A1130609007D
S1131D2893060A0097220000E780C29397220000D6
S1131D38E7800296130405001305040093050400C4
S1131D4897120000E780C26B930A0500374500002C
S1131D589304859D9309000013090000130A600089
S1131D681396F9011305040083A5040063400602D1
S1131D7897120000E780C26893050500130509005F
S1131D8897020000E780C2776F00C0019712000035
S1131D98E7800267930505001305090097220000F0
S1131DA8E780028E1309050093850A0013050400D1
S1131DB897120000E780C264938919001304050090
S1131DC893844400E39E49F98320C1011305090063
S1131DD80324810183244101032901018329C100CA
S1131DE8032A8100832A410013010102678000004D
S1131DF8B706008013C8F6FF130101FF33F8050185
S1131E082326110093880500630E0800B376D500D5
S1131E183707807FB3CEA6001306F7FF6344D601C5
S1131E28635E070197120000E780825D9305050051
S1131E3897120000E780C2B46F00001463CE0E133B
S1131E48638E0E0DB70080001383F0FF634ED30139
S1131E5893958E00930020F8635CB0009380F0FFA4
S1131E68939515006FF05FFF93D57E41938015F825
S1131E78930F20F8634E03011317880013860F008D
S1131E88634C07001306F6FF131717006FF05FFF84
S1131E9813537841130613F863CCF001370E80000E
S1131EA81305FEFFB3FEAE00B3E7CE016F000001D9
S1131EB8930220F8B3831240B3977E00130F20F8DF
S1131EC8634CE601B70F80001388FFFF33F708015E
S1131ED8336FF7016F00C000B308CF40331F1801F8
S1131EE8B388C040B380E741638E08009397170016
S1131EF863C6000063840002939710009388F8FF78
S1131F086FF05FFE63C400009387000063880700D6
S1131F18B7058000938EF5FF6F00000293D2F60197
S1131F28374E000013050EAA93932200B3067500DA
S1131F3803A506006F00400463C8FE0093971700CA
S1131F481306F6FF6FF05FFF130320F86340660281
S1131F58B7028000B3835740130EF607B3E6D300E5
S1131F6813157E0133E5A6006F0000013306C34054
S1131F78B3D7C74033E5D7008320C100130101015B
S1131F886780000093070000638E05001397F5012E
S1131F9863540700B387A70093D5150013151500DC
S1131FA86FF09FFE13850700678000001308050083
S1131FB893030000130500003367D6006302070487
S1131FC89312F60163DC020033030501B338A3005E
S1131FD8B387B30013050300B383F800139EF60117
S1131FE8935EF80113561600139F15003366CE004E
S1131FF893D61600B3E5EE01131818006FF0DFFB53
S1132008938503006780000083254500130101FEC2
S1132018232A910023282101232E1100232C810037
S11320289304050003290500638E05001385050044
S11320382326B10097020000E78082771304050085
S11320486F008001130509002326B10097020000E0
S1132058E7800276130405028325C10013050900ED
S1132068130654FF97020000E78002718320C10120
S113207823A0A4001305C0003305854023A2B4009F
S1132088032481018324410103290101130101026D
S113209867800000130101FB370700802326110421
S11320A89340F7FFB3F315009307F5FF232C41037F
S11320B833B8A7009388F3FF370AF07F232E310340
S11320C8130EFAFFB309180123248104232291046F
S11320D823202105232A510323286103232671037E
S11320E823248103130305001384050093020600C7
S11320F89384060033F91600636E3E036396C901A0
S1132108930AE0FF63E8FA02138BF2FFB33B5B0028
S1132118130CF9FF370FF07FB38E8B01930FFFFF7A
S113212863EADF036394FE0B1307E0FF636467034A
S11321386F00C00963687A00B700F07F639C1300DE
S1132148630A0300370F080093030300B366E4012E
S11321586F00402AB707F07F63E62701631CF90084
S1132168638A02003704080093830200B3E68400FC
S11321786F004028631203026390F3023343940010
S113218863960200B7020080630853321306050001
S1132198938605006F000033639602003708F07FCA
S11321A863020933B3687300B3E92201639A080030
S11321B8639A0930B3735300B37694006F00802395
S11321C81306050093860500638E092E63E6230132
S11321D863107902637E530013050300930504001A
S11321E813830200138404009302050093840500FA
S11321F8B70310001389F3FF1356440193D644011F
S1132208337E2401B3FA24019379F67F13FAF67F17
S113221823286100232AC101232C5100232E5101B4
S1132228639A09001305010197020000E78002DEA2
S113223893090500631A0A00130581019702000037
S1132248E780C2DC130A0500832F41018328C101FA
S1132258832E010103288101370F100033E7EF01B2
S113226833E5E801B3CB8400370B008093D0DE015B
S1132278931737009355D80113133500338A49410E
S11322883379640133FC6B0113943E00B3EBF00023
S1132298B3E46500931A380063180A00232C51012B
S11322A8232E91006F0000069302F00363C44205D5
S11322B8930300043386434113850A00938504007D
S11322C897020000E780424B336EB50013060A00FC
S11322D813850A0093850400333BC001971200005C
S11322E8E78082C5B36EAB00232CD101232EB10045
S11322F86F0040011306100093060000232CC10050
S1132308232ED100032F8101832FC10163060C08FA
S1132318330CE441B33084013387FB41B30B1740DA
S1132328B3677C0123288101232A71011306000065
S11323389306000063880718370480001308F4FF25
S11323486360780B638C0B0013850B0023267101E3
S113235897020000E780C2456F00800113050C0056
S11323682326710197020000E780824413050502C1
S11323788325C100930485FF1386040013050C000C
S113238897020000E780423F2328A100232AB100D6
S1132398B38999406F00C004B308E40133B58800D9
S11323A8B385FB013303B500931A730063C80A00AD
S11323B823281101232A61006F008002131AF301F4
S11323C893D2180033665A0093F3180093561300F7
S11323D8336E76002328C101232AD100938919007A
S11323E8130BE07F635C3B01B70EF07F930300009F
S11323F8B366D901138603006F00C00C6348300527
S1132408032C0101832B41011386F90313050C00E6
S113241893850B0097020000E7800236130F100023
S1132428B36EB50033063F4113050C0093850B00CA
S11324383334D00197120000E78002B0B369A400D6
S113244823283101232AB100930900008320410184
S1132458832F0101139549019397900093D8C700DE
S11324681397D00193D43F003369190113F87F00FF
S113247893054000B3639700B366A90063DE0501C2
S1132488138E1300333B7E00B30BDB0093030E0063
S113249893860B006FF01FF6E31EB8F413F31300D2
S11324A8B38A630033BA7A003306DA0093830A00E6
S11324B8930606006FF01FF437440000032604A3B4
S11324C8832644A38320C1041305060093850600CC
S11324D80324810483244104032901048329C103B7
S11324E8032A8103832A4103032B0103832BC1029B
S11324F8032C81021301010567800000130101FD0B
S113250837070080232611029340F7FFB707807F1F
S1132518B37615009388F6FF1386E7FF232021037B
S1132528232861012324810223229102232E3101CD
S1132538232C4101232A5101232671011309050083
S1132548138B0500B3F2150013880700636816019E
S11325581383F2FF636C66006F00C00563F8D7004D
S1132568370E4000B365C5016F00C01DB703807FF7
S113257863785800370A4000B3654B016F00801C2C
S1132588639C760033496901370B00806308691B33
S1132598930505006F00001B6386721A6398060092
S11325A86392021AB37569016F00C0199305050097
S11325B8638A021863F856001304090013090B0010
S11325C8130B040093547901B7058000938AF5FF2F
S11325D813557B0193F4F40F337A59019379F50F6A
S11325E8B37A5B016390040213050A0097020000A2
S11325F8E780021C930B85FF130E9000331A7A01AF
S1132608B304AE406390090213850A0097020000E0
S1132618E780021A930985FF930E9000B39A3A0152
S1132628B389AE4037078000370F0080B34F2B01C2
S1132638B366EA00B3E8EA0033863441B37BE901C0
S1132648B3F0EF01939236009397380063060602BD
S11326581308F0016340C802930300023384C340A3
S11326683399870033D3C700333B2001B3676B002A
S11326786F00800093071000638C00023384F240DB
S1132688930500006300040C370E0004930AFEFF50
S113269863EE8A021305040097020000E7804211E2
S11326A89309B5FF33143401B38434416F004003F4
S11326B83384570013154400635A050093751400B6
S11326C8135A14003364BA0093841400930EE00F71
S11326D863D89E00B704807FB3E59B006F00800633
S11326E8634290021387F401130F1000B30F9F4045
S11326F8B316E400B350F401B332D00033E412004B
S113270893040000131664001358960093977401F9
S11327183363F800B365730193787400930B400036
S113272863D61B01938515006F00C001639C780173
S113273893F31500B38575006F00C000374500009A
S11327488325C5A38320C1021385050003248102C0
S113275883244102032901028329C101032A810137
S1132768832A4101032B0101832BC10013010103B7
S1132778678000009317A60163D8070013070000B9
S1132788B315C5006F00000263000602930200023D
S11327983383C240B3536500B395C5003317C500EE
S11327A8B3E5B3001305070067800000B707FFFF10
S11327B8B372F50013B31200131743009305000115
S11327C8B383E540B706010033557500138606F058
S11327D83378C50093381800139E3800930E800090
S11327E8338FCE41B35FE50193F20F0F13B3120099
S11327F8B307EE009305400013172300B383E540A5
S113280833D57F009376C50093B8160013082000CB
S1132818139E1800B30EC841335FD5013386E70011
S113282893571F0093C2170013F312003307604035
S1132838B305E841B30FC601B373B70033857F000E
S113284867800000B707008093C2F7FF13070500ED
S113285833F855003705F07F636C05076314A80047
S11328686318070633F35600B703F07F63E2630681
S113287863147300631E0604B70E008033EED5009C
S113288813CFFEFFB368C700B37FEE01B3E7F801C7
S11328981305000063840704B3F2D50063CA020079
S11328A863CCD502639CB600637AC7006F00C0028C
S11328B863C4B6026394D5006360E6023346C70076
S11328C8B3C6D500B365D6003335B00067800000C1
S11328D813051000678000001305F0FF67800000EF
S11328E8370700809342F7FF9307050033F3550039
S11328F83705F07F33F85600636A65066314A3004E
S11329086396070663640507B703F07F63147800CA
S1132918631E0604B70E008033EED50013CFFEFF06
S1132928B3E8C700B37FEE0133E7F80113050000ED
S113293863000704B3F2D50063CA020063C8D50272
S1132948639CB60063FAC7006F00400263C0B60216
S11329586394D500636CF60033C6C700B3C6D500CC
S1132968B365D6003335B000678000001305F0FF67
S11329786780000097020000678002ED130101FDE3
S1132988232C4101135A750123286101137AFA0F84
S1132998370B800023261102232481029300FBFFB6
S11329A8232E3101232671013344B50093DB7501CD
S11329B8B70900801307FAFF9307D00F2322910267
S11329C823202103232A510193FBFB0F3374340181
S11329D8B374150033FB150063E6E7009382FBFF2D
S11329E863FA570A13C3F9FFB3736500B706807F08
S11329F863F8760037034000336565006F004022B2
S1132A0833F9650063F82601370B400033E56501A7
S1132A186F0000216398D300336574006312792032
S1132A286F00801F6302D91C639603006306091EA6
S1132A386F00801B3365D4006304091E37058000CA
S1132A489305F5FF930A000063E0750213850400FB
S1132A5897020000E780C2D5130685FF130890008B
S1132A68B394C400B30AA840B7088000138EF8FFD3
S1132A7863642E0313050B0097020000E78042D31A
S1132A88930E85FF338FAA00331BDB01930A7FFF64
S1132A986F008000930A0000B70F8000B369FB0140
S1132AA8B7F00475330A7A4113873033B30B5A01EC
S1132AB8939A89003309574113860A009306000044
S1132AC81305090093050000B3E4F40197F2FFFF2E
S1132AD8E780024E3305B040130609009306000050
S1132AE89305000097F2FFFFE780824C9397150047
S1132AF89352F50133EB570013860A00930600003E
S1132B0813050B009305000097F2FFFFE780424A84
S1132B183305B04013060B0093060000930500002C
S1132B2897F2FFFFE780C248139315009353F5010A
S1132B38336A730013860A009306000013050A001B
S1132B489305000097F2FFFFE78082463305B04003
S1132B5813060A00930600009305000097F2FFFF8E
S1132B68E7800245939615001355F501B3E5A600D1
S1132B781385E5FF139614009305000093060000DF
S1132B8897F2FFFFE780C242370600011308F6FFF9
S1132B98938A05006362B8021385050093850900CA
S1132BA89394840197F2FFFFE780023EB388A44020
S1132BB8938BFBFF6F00000293DA150013850A005C
S1132BC8938509001399740197F2FFFFE780C23BCC
S1132BD8B308A940138EFB07930EE00FB702807F5A
S1132BE863C8CE036346C001130504006F004003A5
S1132BF8370F8000930FFFFFB3FBFA0193107E0198
S1132C089397180033E77001B3B9F900B302370199
S1132C1833E582006F00C000374400000325C4A3D5
S1132C288320C1020324810283244102032901026F
S1132C388329C101032A8101832A4101032B01014C
S1132C48832BC1001301010367800000130101FFF6
S1132C5823229100B704008093C7F4FF2324810042
S1132C68370780FF3374F500B702007F232611006D
S1132C781383F2FFB300E40023202101B374950009
S1132C88636C1300135734001315D4013704003848
S1132C98330687006F008007B703807F9385F3FFAF
S1132CA863F08502370F4000B377E501930FFFFF08
S1132CB813D837003375F501B70EF07F6F000004A1
S1132CC8630204041305040097020000E78042AE7F
S1132CD813090500930500001305040013065901A0
S1132CE897020000E78042A993089038B7061000BD
S1132CF8338E284133C8B600931E4E0133E60E01C5
S1132D086F00C00013050000130600008320C100F3
S1132D18B36496009385040003248100832441004E
S1132D28032901001301010167800000935775010D
S1132D383707800093F2F70F9305F7FF9356F54191
S1132D483373B500130101FF138612F813056001EC
S1132D5823261100B363E30093E01600636CC500F7
S1132D6893087001338EC84013850000B3D5C3019E
S1132D786F00800113050000634C06001388A2F657
S1132D8813850000B395030197F2FFFFE780C21F84
S1132D988320C100130101016780000013567501E7
S1132DA89372F60F938512F81308000063CA05029C
S1132DB863480502B70680009387F6FF3373F5006E
S1132DC8930370013367D30063D8B3009388A2F6E2
S1132DD8331817016F00C0003385B3403358A70078
S1132DE81305080067800000130101FF23248100F4
S1132DF82326110023229100232021011304050016
S1132E08630E050493040000635605003304A040D0
S1132E18B70400801305040097020000E780429974
S1132E281309050013065901130504009355F441C9
S1132E3897020000E78042949307E04137071000A7
S1132E48B3822741B3C5E50013934201B303B3002A
S1132E5833E69300930506006F00C00013050000D5
S1132E68930500008320C1000324810083244100CA
S1132E78032901001301010167800000130101FF08
S1132E882324810013040500232611002322910022
S1132E981305000063060408930400006356040045
S1132EA833048040B704008013050400970200002F
S1132EB8E78002901307F001B302A740930670015C
S1132EC8B707800063CA5600930E85FF331FD401E9
S1132ED8334EFF006F008003930080003383A040CB
S1132EE893058501B35364003316B4003708008092
S1132EF833CEF3006376C800130E1E006F00000182
S1132F086316060193781E00330E1E01930FE00921
S1132F183385AF401314750133078E00336597006A
S1132F288320C1000324810083244100130101018B
S1132F38678000009317A60163D8070013070000F1
S1132F4833D5C5006F000002630006029302000235
S1132F583383C24033D7C500B39365003356C500E5
S1132F6833E5C30093050700678000008325450007
S1132F78130101FE232A910023282101232E110085
S1132F88232C81009304050003290500638E0500A2
S1132F98138505002326B10097020000E7804281CB
S1132FA8130405006F008001130509002326B100EE
S1132FB897F2FFFFE780C27F130405028325C1004F
S1132FC813050900130654FF97F2FFFFE780C27A3E
S1132FD88320C10123A0A4001305C0003305854044
S1132FE823A2B4000324810183244101032901019C
S1132FF81301010267800000130101FA13D7450188
S1133008B70210001383F2FF23244105137AF77FD4
S1133018232E1104232821052326310593D04601A4
S1133028B3C7D50037090080B3F3650033F86600E9
S11330389308FAFF9309D07F232C8104232A91044F
S11330482322510523206105232E7103232C810398
S1133058232A91032328A1032326B10393FAF07F9B
S113306813040000B3F427012328A100232A7100C4
S1133078232CC100232E010163E61901138BFAFFE7
S113308863F8690D934BF9FF33FB7501370CF07F37
S113309863666C01631C8B01630A0500B7060800AC
S11330A893020500B3E0D5006F000030B3FC76014D
S11330B8B705F07F63E69501639CBC00630A0600CC
S11330C8B708080013050600B3E516016F00402F82
S11330D8631C0500631ABB003365960113080400DA
S11330E8631A051A6F00002DB366650163100602A2
S11330F8B70DF07F639CBC01638E062A33EE9401FE
S11331081305040093050E006F00802B6386061ACE
S1133118336F960163020F1AB70F10001389FFFF6C
S1133128130D0000636A6901130501019702000089
S1133138E78002E4130D0500636E9901130581010C
S113314897020000E780C2E2330DAD006F008000F3
S1133158130D0000832781010327C101832901017D
S113316883204101B70B1000B3627701139CB700A9
S113317813D357019393B2001386090013050C0067
S11331889306000093050000B36C73002326110016
S113319897F2FFFFE780C2E1138B0500138609004D
S11331A8930D05009306000013850C009305000099
S11331B897F2FFFFE780C2DF0328C1001309050067
S11331C893890500B36878011386080013050C0079
S11331D893060000930500002326110197F2FFFFD0
S11331E8E78002DDB3066901032EC100338BA60014
S11331F833B626013335DB00338C35013309C5007A
S11332089305000013850C0013060E0093060000B6
S113321897F2FFFFE780C2D9B30EAC00B3393C0183
S1133228B385B900B3872E0133BF8E01B30FBF0036
S113323833B7D701B309F701938A1AC0338A4A010D
S11332489392B900938B0D00938C0700330DAA0158
S113325863D60200130D1D006F00C002939B190072
S11332689353FB0193D0F7011393170013D8FD016F
S1133278131B1B00B3E97001B3EC6300939B1D009F
S1133288336B6801930DE07F63DEAD01130804001E
S1133298370BF07FB3EB64011305080093850B002B
S11332A86F000012634EA009130C1000330AAC41DE
S11332B8130EF00363584E011305040093850400AC
S11332C86F00001013850B0093050B0013060A000A
S11332D897020000E78042C6130DFD03930D050015
S11332E8938A050013060D0013850C0093850900C5
S11332F897F2FFFFE780424833E9AD0033ECBA00A8
S113330813850B0093050B0013060D0097F2FFFFBE
S1133318E7808246B36EB500333FD00113850C00B5
S11333289385090013060A00B36BE90197020000AC
S1133338E78082C0130B0C00130905006F00C0015D
S1133348B70810009386F8FF33F6D90013154D011A
S113335813890C00B365C500B36289003704008083
S1133368B3E095006366640163108B0263800B020B
S113337813831200B3335300B38913009302030079
S1133388938009006F00400263900B02631E8B0058
S113339893F41200B3859200B3BF5500B3871F009E
S11333A8938205009380070013850200938500002B
S11333B86F000001B74E000003A50EA383A54EA31A
S11333C88320C105032481058324410503290105BC
S11333D88329C104032A8104832A4104032B010499
S11333E8832BC103032C8103832C4103032D010385
S11333F8832DC1021301010667800000130101FE39
S1133408232A910093547501232631012322510163
S1133418B709800093FAF40F9382F9FF232E110061
S1133428232C81002328210193D075013344B5004E
S1133438370900801387FAFF9307D00F232061010F
S11334482324410193F4F00F33742401337B550092
S1133458B3F9550063E6E7001383F4FF63FE670AD4
S11334689343F9FF33767500B706807F63F8C60087
S1133478B7084000336515016F00001C33F9750067
S113348863F82601370B400033E565016F00C01A65
S11334986318D6003365C4006310091A6F00401915
S11334A86318D90033652401631806186F0040189F
S11334B86304060063160900130504006F00C017AF
S11334C8370580009305F5FF130A000063E0C50281
S11334D813050B0097F2FFFFE780822D130885FF81
S11334E893089000331B0B01338AA840370E8000E1
S11334F8930EFEFF63E42E031385090097F2FFFF82
S1133508E780022B130F85FFB30FAA40B399E90193
S1133518138A9F006F008000130A0000B700800020
S1133528B3E21900139582009305000033661B006B
S11335389306000097F2FFFFE78082A7938414F8AC
S1133548B38A540113938500938305001309050076
S1133558B3874A0163560300938717006F0040013D
S1133568139A15001357F501B363EA0013191500EC
S11335781306E00F6358F600B705807F3365B4007F
S11335886F00800B634AF00693081000338EF840EE
S1133598930EF00163C4CE03338AD7013357C901AC
S11335A83396430133194901B366C7003335200103
S11335B833E9A60033DBC3016F004005130FF003A2
S11335C86344CF03B38FE701B390F301930A10FE6A
S11335D8B3E22001B387FA40B334500033D3F30085
S11335E833E964006F00C000B3E9230133393001C3
S11335F8130B00006F008001B70680001385F6FFE7
S1133608B3F5A30013987701336BB80033658B00C7
S11336183704008063762401130515006F00C00188
S1133628631C890093731500330575006F00C0008F
S1133638374800000325C8A38320C101032481015E
S113364883244101032901018329C100032A81003C
S1133658832A4100032B0100130101026780000043
S11336681307060037060080B3C7C6009386070011
S11336781306070097F2FFFF678002A2B7070080CE
S1133688B3C5F50097F2FFFF678082E7130101FED7
S1133698232A9100B704008013C6F4FF232E1100D7
S11336A8370710B8B3F0C500B707F0C7B382E00016
S11336B83383F000232C81002328210123263101A0
S11336C82324410113040500B3F4950063685300EF
S11336D8B703F07F63F213046F008004B706002079
S11336E89388F6FF139530001358D401B375140169
S11336F8B7090010336A05013709004063F8B900B7
S1133708930E1900B302DA016F00800DB3022A0187
S11337186398350D6F00C00B63907002630E05004B
S1133728B70040009387F0FF3373F400B703C07FFA
S1133738B36273006F00C00A3705F0476360150A67
S11337486394A000631C040813D84001130A1038BA
S1133758330A0A41930640039302000063C24609F0
S1133768B70810009389F8FFB3F53501B3E91501DB
S11337781306F8CB130504009385090097F2FFFF9D
S1133788E78082FF3369B50013060A0013050400B5
S11337989385090097F2FFFFE780027A3339200105
S11337A8B70F0020336EA9001384FFFF939E3500E2
S11337B8135FDE0133768E0037070010B3E2EE01A3
S11337C86376C700938212006F008001631AE600D3
S11337D813FE1200B382C2016F008000B702807F1B
S11337E88320C10133E5920003248101832441012C
S11337F8032901018329C100032A8100130101025D
S107380867800000D1
S11338100000404000002041000040410000C04042
S11338200000A040000000420000003F0000803F74
S113383000005842000000400000804000000000EA
S11338409A9999999999D93F9A9999999999E93F06
S1133850343333333333F33F9A9999999999F93F30
S1133860000000000000004034333333333303409E
S113387067666666666606409A99999999990940B9
S1133880CDCCCCCCCCCC0C400000000000001040CF
S11338909A999999999911403433333333331340B6
S11338A09A9999999999B93FF0F89C8E8783878E54
S11338B09CF8F00000FEFF0303030303070EFCF86B
S11338C00000FEFF0303030303070EFCF80000FFE0
S11338D0FF00000000000000FFFF0000FEFF8383E4
S11338E0838383C7EE7C380000F8FC0E07030303D0
S11338F0070EFCF800003F7FE0C08080C0E07F3FFF
S1133900FFFF01010101010101FFFF0000FFFF0CA6
S11339100C0C0C1C3E77E3C100007FFFC0C0C0C08C
S1133920C0E0703F1F00001F3F70E0C0C0C0E070E7
S11339303F1F00007FFFC1C1C1C1C1E3773E1C002E
S1133940001F3F70E0C0C0C0E0703F1F00000000D7
S11339500001FFFF0100000000FF00FF00FF00FF67
S113396000FF00FF00FF00FF00FF00FF00FF00FF5B
S113397000FF5AFF00FF00FF00FF00FF00FF00FFF1
S113398000FF00FF00FF00FF00FF00FF00FF00FF3B
S113399000FF00FF00FF00FF03FF0BFF13FF1BFFEF
S11339A023FF2BFF33FF3BFF43FF4BFF53FF5BFF23
S11339B063FF6BFF73FF7BFF83FF8BFF93FF9BFF13
S11339C0A3FFABFFB3FFBBFFC3FFCBFFD3FFDBFF03
S11339D0E3FFEBFFF3FFFBFF0000803FABAA2A3EAF
S11339E08988083C010D50391DEF38362B32D73207
S10739F05804000073
S11339F40000000000FFFFFF10FFFFFF00F8FFFFBF
S1133A08182D4454FB210940182D4454FB21194016
S1133A18182D4454FB2109C0182D4454FB21F93FA7
S1133A28182D4454FB21F9BF000000000000F87F62
S1133A38DB0FC9400000C07F000000000000000048
S1133A48F8FE373337FEF800FFFFC9C9C9FF76000F
S1133A58FFFFC1C1C1FF7E00FFFFDBDBDBC3C30087
S1133A68FFFF181818FFFF00FFFFC0C0C0C0C00048
S1133A78FFFFC3C3C3FFFF00FFFF090919FFF600D7
S1133A887FFFC0C0C0FF7F000F1FD8D8D8FFFF003A
S1133A988100000080000000000000000000008099
S9030400F8
                                                                                                                                                                                                                                                                                                                                       